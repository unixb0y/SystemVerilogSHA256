`default_nettype none
`timescale 1 ns / 10 ps

module sha_mainloop_tb;
	logic [511:0] padded;
	logic clk, rst;

	sha_mainloop uut(.padded(padded), .clk(clk), .rst(rst));

	initial begin
    	$dumpfile("sha_mainloop_tb.vcd");
    	$dumpvars;
    	assign padded = 512'b01100001011000100110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000;
    	assign clk = 0;
    	assign rst = 1;
    	#5;
    	assign clk = 1; #5
    	assign rst = 0; #5
    	for(int i=0; i<150; i++) begin
    		assign clk = ~clk;
    		#5;
    	end
    	$display("FINISHED mainloop_tb");
    	$finish;
	end
endmodule